grammar concretesyntax;

imports abstractsyntax;
synthesized attribute unparse :: String;
