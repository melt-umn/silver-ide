grammar parsers;

import concretesyntax as cst;
import concretesyntax:regex;
import silver:definition:regex;

parser specFileParser :: cst:SpecRoot {
  concretesyntax;
  concretesyntax:regex;
  silver:definition:regex;
}
