grammar parsers;

imports concretesyntax as cst;

parser specFileParser :: cst:SpecRoot {
  concretesyntax;
}
