grammar parsers;

import concretesyntax:specList;

parser specNameListParser :: SpecNameList {
  concretesyntax:specList;
}
