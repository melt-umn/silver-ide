grammar slide:parsers;

imports slide:concretesyntax as cst;

parser specFileParser :: cst:SpecRoot {
  slide:concretesyntax;
}
