grammar abstractsyntax;

{-- attributes occuring on terminals, nonterminals and lexer classes --}
synthesized attribute atomMarkupName:: Maybe<String>;
