grammar slide:concretesyntax;

imports slide:abstractsyntax;
synthesized attribute unparse :: String;
